module ALUControl (
    input [1:0] ALUOp,
    input [5:0] funct,
    output reg [3:0] alu_control
);
always @(*) begin
    case (param)
        : 
        default: 
    endcase
end
    
endmodule